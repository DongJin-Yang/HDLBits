module top_module ( input a, input b, output out );
    mod_a instance_1(a, b, out);
endmodule

